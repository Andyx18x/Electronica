module comp_and(input wire a, 
                input wire b,
                output wire x);

assign x = a & b;

endmodule
